module VGA_top(
input CLK,
input RX,
output TX,
output VGA_HS, VGA_VS, 
output VGA_R0, VGA_R1, VGA_R2, 
output VGA_G0, VGA_G1, VGA_G2, 
output VGA_B0, VGA_B1, VGA_B2,
output S1_A, S1_B, S1_C, S1_D, S1_E, S1_F, S1_G,
output S2_A, S2_B, S2_C, S2_D,S2_E, S2_F, S2_G);


